library verilog;
use verilog.vl_types.all;
entity tb_obp is
end tb_obp;
