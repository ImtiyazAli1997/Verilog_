library verilog;
use verilog.vl_types.all;
entity tb_exor is
end tb_exor;
