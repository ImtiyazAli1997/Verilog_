library verilog;
use verilog.vl_types.all;
entity hw1 is
    port(
        y1              : out    vl_logic;
        y0              : out    vl_logic;
        i               : in     vl_logic;
        s               : in     vl_logic
    );
end hw1;
