library verilog;
use verilog.vl_types.all;
entity basic_gates_tb is
end basic_gates_tb;
