library verilog;
use verilog.vl_types.all;
entity my_not_tb is
end my_not_tb;
