library verilog;
use verilog.vl_types.all;
entity sub is
end sub;
