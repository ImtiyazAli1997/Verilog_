module my_not(
	input a,
	output y);
	
	not n1 (y,a);
	
endmodule