module mul8_v2 (input [7:0] a,b, output [15:0] y);

	genvar i,j;
	wire [7:0]p[0:7];
	//wire [7:0] p[0];
	//wire [7:0] p[1]
	//wire [7:0] p[2]
	//wire [7:0] p[3]
	//wire [7:0] p[4]..
	
	
	//the block outside the alwaus is generator block
	
	for(i=0;i<8;i=i+1)	begin
		for (j=0;j<8;j=j+1) begin
			and Gij	(p[i][j],a[i],b[j]);
		end
	end
	
	
	wire [14:0] R0,R1,R2,R3,R4,R5,R6,R7;
	
	assign R0 = {7'b0000000,p[0][7],p[0][6],p[0][5],p[0][4],p[0][3],p[0][2],p[0][1],p[0][0]};
	assign R1 = {6'b000000,p[1][7],p[1][6],p[1][5],p[1][4],p[1][3],p[1][2],p[1][1],p[1][0],1'b0};
	assign R2 = {5'b00000,p[2][7],p[2][6],p[2][5],p[2][4],p[2][3],p[2][2],p[2][1],p[2][0],2'b00};
	assign R3 = {4'b0000,p[3][7],p[3][6],p[3][5],p[3][4],p[3][3],p[3][2],p[3][1],p[3][0],3'b00};
	assign R4 = {3'b00,p[4][7],p[4][6],p[4][5],p[4][4],p[4][3],p[4][2],p[4][1],p[4][0],4'b0000};
	assign R5 = {2'b00,p[5][7],p[5][6],p[5][5],p[5][4],p[5][3],p[5][2],p[5][1],p[5][0],5'b00000};
	assign R6 = {1'b0,p[6][7],p[6][6],p[6][5],p[6][4],p[6][3],p[6][2],p[6][1],p[6][0],6'b000000};
	assign R7 = {p[7][7],p[7][6],p[7][5],p[7][4],p[7][3],p[7][2],p[7][1],p[7][0],7'b0000000};
	
	assign y=R0+R1+R2+R3+R4+R5+R6+R7;
endmodule
			