library verilog;
use verilog.vl_types.all;
entity tb_nand is
end tb_nand;
