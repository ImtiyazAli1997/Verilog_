library verilog;
use verilog.vl_types.all;
entity tb_and is
end tb_and;
