library verilog;
use verilog.vl_types.all;
entity tb_not is
end tb_not;
