library verilog;
use verilog.vl_types.all;
entity tb4 is
end tb4;
