library verilog;
use verilog.vl_types.all;
entity tb_or is
end tb_or;
